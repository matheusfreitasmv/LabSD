-- Questão 2 letra (a)

library  ieee;
use ieee.std_logic_1164.all;

entity ex_2 is
